LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.All;

ENTITY mips is --single cycle MIPS processor
	PORT(
		clk, reset: IN STD_LOGIC;
		pc: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		instr: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		memwrite: OUT STD_LOGIC;
		aluout, writedata: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		readdata: IN STD_LOGIC_VECTOR(31 DOWNTO 0));
END mips;

Architecture Behavioral of mips IS

	--Universal
	SIGNAL INSTRUCTION_TYPE: STD_LOGIC;
	SIGNAL REGISTER_SOURCE_ADDRESS: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL REGISTER_DESTINATION_ADDRESS: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL FUNCTION_CODE: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL REGISTER_TEMP_ADDRESS: STD_LOGIC_VECTOR(5 DOWNTO 0);
	--R Type
	SIGNAL R_IMMEDIATE_VALUE: STD_LOGIC_VECTOR(8 DOWNTO 0);
	--I Type
	SIGNAL I_IMMEDIATE_VALUE: STD_LOGIC_VECTOR(14 DOWNTO 0);
	
	BEGIN
		INSTRUCTION_TYPE <= instr(0)
		REGISTER_SOURCE_ADDRESS <= instr(6 DOWNTO 1);
		REGISTER_DESTINATION_ADDRESS <= instr(12 DOWNTO 7);
		FUNCTION_CODE <= instr(16 DOWNTO 13);
		IF (INSTRUCTION_TYPE='0') THEN--R Type
			REGISTER_TEMP_ADDRESS <= instr(22 DOWNTO 17);
			R_IMMEDIATE_VALUE <= instr(31 DOWNTO 23);
		ELSIF (INSTRUCTION_TYPE='1') THEN--I Type
			I_IMMEDIATE_VALUE <= instr(31 DOWNTO 17);
		END IF;
		
END Behavioral;
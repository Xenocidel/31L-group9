LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.All;

PACKAGE comp_pkg IS
	--mips--
	
	--alu--
	
	--dma--
	
	--instruction memory (cache)--
	
	--pc--
	
	--sign extender--
	
	--regfile--
	
	--mux--
	
END comp_pkg;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.All;

ENTITY fifo IS
	GENERIC(NBIT : INTEGER := 32;
			DEPTH : INTEGER := 4);
	PORT (

		);
END fifo ;

ARCHITECTURE Structural OF fifo IS
	
	BEGIN
	
END Structural;
module mips_tb ();

	bit clk, clk_mips, rst, req, ack;
	logic [5:0] dma_addr, dma_addrout, instr_addr;
	logic [31:0] dma_data, dma_dataout, instr_data;
	reg [31:0] main_mem [63 :0];
	logic [31: 0] data_out, instruction, instruct_out; 
	integer x; 
	
	dma D1(
        .clk(clk)
        ,.rst(rst)
        ,.req(req)
        ,.addr(dma_addr)
        ,.data(dma_data)
        ,.ack(ack)
		,.addr_o(dma_addrout)
		,.data_o(dma_dataout)
        );
	
	controllermips C1(
		.clk(clk)
		,.reset(rst)
		,.addr(instr_addr)
		,.instruction(instruction)
		,.data_out(data_out)
		,.instruct_out(instruct_out)
	);
	initial begin 
	
	clk = 1'b0;
	rst = 1'b1; 
	//Main Memory (64 addresses)
	main_mem [0] <= 32'b10000000000011011111111111111111;
	main_mem [1] <= 32'b10000010000101011011111111111101;
	main_mem [2] <= 32'b10000100000111011000000110111111;
	main_mem [3] <= 32'b10000110001001011101101010001001;
	main_mem [4] <= 32'b00000010001010000000010000000000;
	main_mem [5] <= 32'b00000100001100001000011000000000;
	main_mem [6] <= 32'b00001000001110010000010000000000;
	main_mem [7] <= 32'b00000010010000011000100000000000;
	main_mem [8] <= 32'b00001000010010101000011000000000;
	main_mem [9] <= 32'b00000110010100110000001000000000;
	main_mem [10] <= 32'b00000010010110111000010000000000;
	main_mem [11] <= 32'b00000010011001000000100000000000;
	main_mem [12] <= 32'b00000100011011001000001000000000;
	main_mem [13] <= 32'b00001000011101011000010000000000;
	main_mem [14] <= 32'b00000110011111011000100000000000;
	main_mem [15] <= 32'b00000100100001001000011000000000;
	main_mem [16] <= 32'b00001000100011000000001000000000;
	main_mem [17] <= 32'b00000010100100111000010000000000;
	main_mem [18] <= 32'b00000100100110110000100000000000;
	main_mem [19] <= 32'b00001000101000101000001000000000;
	main_mem [20] <= 32'b00000110101010011000010000000000;
	main_mem [21] <= 32'b00000100101100010000100000000000;
	main_mem [22] <= 32'b00001000101110001000001000000000;
	main_mem [23] <= 32'b00000110110000000000010000000000;
	main_mem [24] <= 32'b00000010110010000000100000000000;
	main_mem [25] <= 32'b00001000110100001000001000000000;
	main_mem [26] <= 32'b00000110110110010000010000000000;
	main_mem [27] <= 32'b00000100111000011000100000000000;
	main_mem [28] <= 32'b00000110111010101000001000000000;
	main_mem [29] <= 32'b00000110111100110000100000000000;
	main_mem [30] <= 32'b00000010111110111000010000000000;
	main_mem [31] <= 32'b00001001000001000000001000000000;
	main_mem [32] <= 32'b00000011000011011000010000001011;
	main_mem [33] <= 32'b00001001000101011000100000001011;
	main_mem [34] <= 32'b00000111000111011001000000001011;
	main_mem [35] <= 32'b00000101001001011001011000001111;
	main_mem [36] <= 32'b10000101001010000001001000010000;
	main_mem [37] <= 32'b10001001001100001000101000000000;
	main_mem [38] <= 32'b10000011001110010001001000000000;
	main_mem [39] <= 32'b10001001010000011010010000000000;
	main_mem [40] <= 32'b10000111010010101001011000000000;
	main_mem [41] <= 32'b10000011010100110010010000000000;
	main_mem [42] <= 32'b10000011010110111100100000000000;
	main_mem [43] <= 32'b10000101011001000100100000000000;
	main_mem [44] <= 32'b10001001011011001100101000000000;
	main_mem [45] <= 32'b10000111011101011100110000000000;
	main_mem [46] <= 32'b10000101011111011110110000000000;
	main_mem [47] <= 32'b10001001100001001010110000000000;
	main_mem [48] <= 32'b10000011100011000011101000000000;
	main_mem [49] <= 32'b10001001100100111000001000000000;
	main_mem [50] <= 32'b10000011100110110000000000000000;
	main_mem [51] <= 32'b10000101101000101000100000000000;
	main_mem [52] <= 32'b10001001101010011000001000000000;
	main_mem [53] <= 32'b10000111101100010000100000000000;
	main_mem [54] <= 32'b10000101101110001000110000000000;
	main_mem [55] <= 32'b10001001110000000000111000000000;
	main_mem [56] <= 32'b10000111110010001001000000000000;
	main_mem [57] <= 32'b10000011110100010001001000000000;
	main_mem [58] <= 32'b10000101101110011010000000000000;
	main_mem [59] <= 32'b10000101111000101100010000000000;
	main_mem [60] <= 32'b10000011111010110000010000000000;
	main_mem [61] <= 32'b10001001111100111000001000000000;
	main_mem [62] <= 32'b10000111111111000000000000000000;
	main_mem [63] <= 32'b10000010000000000000000000000000;
	
	for (x = 0; x < 64; x = x + 1) begin		//Load instructions from main memory through DMA to instruction memory
		#50;
		instruction = main_mem[x];
		instr_addr = x;
		$display("Main Memory: Instruction %b \n address: %d", instruction, instr_addr); 
		#50;
	end
	rst = 1'b0;
	#50000;
	
	$finish;
end

always #50 clk = ~clk;

always @ (posedge clk) begin
	if (rst == 0) begin
		$display("\n Data Out: %b", data_out);
		$display("\n Instruct Out: %b", instruct_out); 
	end
end

		
		

endmodule	
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity encoder IS
	PORT(
	in0:IN std_logic;
	in1:IN std_logic;
	f:OUT std_logic;
	);
end encoder;

architecture lab1 of encoder IS
begin
	f <= ;
end lab1;